//----------------------------------------------------------------------
// Created with uvmf_gen version 2023.4_2
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//     
// DESCRIPTION: This file contains macros used with the fsm_out package.
//   These macros include packed struct definitions.  These structs are
//   used to pass data between classes, hvl, and BFM's, hdl.  Use of 
//   structs are more efficient and simpler to modify.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//

// ****************************************************************************
// When changing the contents of this struct, be sure to update the to_struct
//      and from_struct methods defined in the macros below that are used in  
//      the fsm_out_configuration class.
//
  `define fsm_out_CONFIGURATION_STRUCT \
typedef struct packed  { \
     uvmf_active_passive_t active_passive; \
     uvmf_initiator_responder_t initiator_responder; \
     } fsm_out_configuration_s;

  `define fsm_out_CONFIGURATION_TO_STRUCT_FUNCTION \
  virtual function fsm_out_configuration_s to_struct();\
    fsm_out_configuration_struct = \
       {\
       this.active_passive,\
       this.initiator_responder\
       };\
    return ( fsm_out_configuration_struct );\
  endfunction

  `define fsm_out_CONFIGURATION_FROM_STRUCT_FUNCTION \
  virtual function void from_struct(fsm_out_configuration_s fsm_out_configuration_struct);\
      {\
      this.active_passive,\
      this.initiator_responder  \
      } = fsm_out_configuration_struct;\
  endfunction

// ****************************************************************************
// When changing the contents of this struct, be sure to update the to_monitor_struct
//      and from_monitor_struct methods of the fsm_out_transaction class.
//
  `define fsm_out_MONITOR_STRUCT typedef struct packed  { \
  bit _idle_o ; \
  bit _auto_zero_o ; \
  bit _integrate_o ; \
  bit _deintegrate_o ; \
  bit _ref_sign_o ; \
  bit _interrupt_o ; \
  bit [11:0] _measurement_count_o ; \
     } fsm_out_monitor_s;

  `define fsm_out_TO_MONITOR_STRUCT_FUNCTION \
  virtual function fsm_out_monitor_s to_monitor_struct();\
    fsm_out_monitor_struct = \
            { \
            this._idle_o , \
            this._auto_zero_o , \
            this._integrate_o , \
            this._deintegrate_o , \
            this._ref_sign_o , \
            this._interrupt_o , \
            this._measurement_count_o  \
            };\
    return ( fsm_out_monitor_struct);\
  endfunction\

  `define fsm_out_FROM_MONITOR_STRUCT_FUNCTION \
  virtual function void from_monitor_struct(fsm_out_monitor_s fsm_out_monitor_struct);\
            {\
            this._idle_o , \
            this._auto_zero_o , \
            this._integrate_o , \
            this._deintegrate_o , \
            this._ref_sign_o , \
            this._interrupt_o , \
            this._measurement_count_o  \
            } = fsm_out_monitor_struct;\
  endfunction

// ****************************************************************************
// When changing the contents of this struct, be sure to update the to_initiator_struct
//      and from_initiator_struct methods of the fsm_out_transaction class.
//      Also update the comments in the driver BFM.
//
  `define fsm_out_INITIATOR_STRUCT typedef struct packed  { \
  bit _idle_o ; \
  bit _auto_zero_o ; \
  bit _integrate_o ; \
  bit _deintegrate_o ; \
  bit _ref_sign_o ; \
  bit _interrupt_o ; \
  bit [11:0] _measurement_count_o ; \
     } fsm_out_initiator_s;

  `define fsm_out_TO_INITIATOR_STRUCT_FUNCTION \
  virtual function fsm_out_initiator_s to_initiator_struct();\
    fsm_out_initiator_struct = \
           {\
           this._idle_o , \
           this._auto_zero_o , \
           this._integrate_o , \
           this._deintegrate_o , \
           this._ref_sign_o , \
           this._interrupt_o , \
           this._measurement_count_o  \
           };\
    return ( fsm_out_initiator_struct);\
  endfunction

  `define fsm_out_FROM_INITIATOR_STRUCT_FUNCTION \
  virtual function void from_initiator_struct(fsm_out_initiator_s fsm_out_initiator_struct);\
           {\
           this._idle_o , \
           this._auto_zero_o , \
           this._integrate_o , \
           this._deintegrate_o , \
           this._ref_sign_o , \
           this._interrupt_o , \
           this._measurement_count_o  \
           } = fsm_out_initiator_struct;\
  endfunction

// ****************************************************************************
// When changing the contents of this struct, be sure to update the to_responder_struct
//      and from_responder_struct methods of the fsm_out_transaction class.
//      Also update the comments in the driver BFM.
//
  `define fsm_out_RESPONDER_STRUCT typedef struct packed  { \
  bit _idle_o ; \
  bit _auto_zero_o ; \
  bit _integrate_o ; \
  bit _deintegrate_o ; \
  bit _ref_sign_o ; \
  bit _interrupt_o ; \
  bit [11:0] _measurement_count_o ; \
     } fsm_out_responder_s;

  `define fsm_out_TO_RESPONDER_STRUCT_FUNCTION \
  virtual function fsm_out_responder_s to_responder_struct();\
    fsm_out_responder_struct = \
           {\
           this._idle_o , \
           this._auto_zero_o , \
           this._integrate_o , \
           this._deintegrate_o , \
           this._ref_sign_o , \
           this._interrupt_o , \
           this._measurement_count_o  \
           };\
    return ( fsm_out_responder_struct);\
  endfunction

  `define fsm_out_FROM_RESPONDER_STRUCT_FUNCTION \
  virtual function void from_responder_struct(fsm_out_responder_s fsm_out_responder_struct);\
           {\
           this._idle_o , \
           this._auto_zero_o , \
           this._integrate_o , \
           this._deintegrate_o , \
           this._ref_sign_o , \
           this._interrupt_o , \
           this._measurement_count_o  \
           } = fsm_out_responder_struct;\
  endfunction
// pragma uvmf custom additional begin
// pragma uvmf custom additional end
